library ieee;
USE ieee.std_logic_1164.all; 

entity sipoTb is
end sipoTb;

architecture sipoTb_rtl of sipoTb is
  component SerialInParallelOut is
    port
    (
      clk         : in std_logic;        
      nrst        : in std_logic;        
      SerialIn    : in std_logic;            
      ParallelOut : out std_logic_vector(255 downto 0)
    );    
  end component;

  signal halfClk : time := 10 ns;
  signal fullClk : time := 20 ns;
  signal clk : std_logic := '0';
  signal nrst        : std_logic;        
  signal SerialIn    : std_logic;            
  signal ParallelOut : std_logic_vector(255 downto 0);

  begin
    sipoPortMap : SerialInParallelOut port map
    (
        clk => clk,
        nrst => nrst,
        SerialIn => SerialIn,
        ParallelOut => ParallelOut
    );

    clock : process
      begin
        clk <= not clk;
        wait for halfClk;
      end process;

    test : process
      begin
        report "Test start";
        nrst <= '0';
        wait for halfClk;
        nrst <= '1';
        SerialIn <= '0';
        wait for fullClk;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0110000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1100100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1001011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0111010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1110100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1001111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0011110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1010001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0100010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0101101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1101000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1010001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0010000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0100001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1000011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0000110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0001100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0011000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0110000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1100001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1000010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0000101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"0001011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0010111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011010" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0101110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000110100" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1011101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001101000" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011010000" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000110100001" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1101111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001101000010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1011111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011010000101" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"0111111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000110100001010" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001101000010101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011010000101011" report "sipo has the wrong output" severity failure;
        SerialIn <= '0';
        wait for fullClk;
        assert ParallelOut = b"1111100011101000111001101010111011101111101010100100110110101010100111010101100100111100001100111100011110110010010000000110111001011111101110000000100110000010011001000110011110010101110110000101110010101001101110001110010100110101011101000110100001010110" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1111000111010001110011010101110111011111010101001001101101010101001110101011001001111000011001111000111101100100100000001101110010111111011100000001001100000100110010001100111100101011101100001011100101010011011100011100101001101010111010001101000010101101" report "sipo has the wrong output" severity failure;
        SerialIn <= '1';
        wait for fullClk;
        assert ParallelOut = b"1110001110100011100110101011101110111110101010010011011010101010011101010110010011110000110011110001111011001001000000011011100101111110111000000010011000001001100100011001111001010111011000010111001010100110111000111001010011010101110100011010000101011011" report "sipo has the wrong output" severity failure;
                
      end process;
end sipoTb_rtl;