LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity Testbench is
end Testbench;

architecture tb of Testbench is
  component SBox
    port
    (
      data_in : in std_logic_vector(127 downto 0);
      data_out : out std_logic_vector(127 downto 0)
    );
  end component;

  signal data_in : std_logic_vector(127 downto 0);
  signal data_out : std_logic_Vector(127 downto 0);

  begin
    SBoxPort : SBox port map
    (
        data_in => data_in,
        data_out => data_out
    );

    test : process

    impure function test(data : std_logic_vector(127 downto 0)) return boolean is
      begin
        data_in <= data;
        return true;
    end test;

    impure function as(data : std_logic_vector(127 downto 0)) return boolean is
      begin
        assert data_out = data report "SBox wrong" severity error;
        return true;
    end as;

      variable foo : boolean := false;
      variable delay : time := 2 ns;

      begin
        foo := test(x"00000000000000000000000000000000");
        wait for delay;
        foo := as(x"63636363636363636363636363636363");
        foo := test(x"00000000000000000000000000000001");
        wait for delay;
        foo := as(x"6363636363636363636363636363637C");
        foo := test(x"00000000000000000000000000000002");
        wait for delay;
        foo := as(x"63636363636363636363636363636377");
        foo := test(x"00000000000000000000000000000003");
        wait for delay;
        foo := as(x"6363636363636363636363636363637B");
        foo := test(x"00000000000000000000000000000004");
        wait for delay;
        foo := as(x"636363636363636363636363636363F2");
        foo := test(x"00000000000000000000000000000005");
        wait for delay;
        foo := as(x"6363636363636363636363636363636B");
        foo := test(x"00000000000000000000000000000006");
        wait for delay;
        foo := as(x"6363636363636363636363636363636F");
        foo := test(x"00000000000000000000000000000007");
        wait for delay;
        foo := as(x"636363636363636363636363636363C5");
        foo := test(x"00000000000000000000000000000008");
        wait for delay;
        foo := as(x"63636363636363636363636363636330");
        foo := test(x"00000000000000000000000000000009");
        wait for delay;
        foo := as(x"63636363636363636363636363636301");
        foo := test(x"0000000000000000000000000000000A");
        wait for delay;
        foo := as(x"63636363636363636363636363636367");
        foo := test(x"0000000000000000000000000000000B");
        wait for delay;
        foo := as(x"6363636363636363636363636363632B");
        foo := test(x"0000000000000000000000000000000C");
        wait for delay;
        foo := as(x"636363636363636363636363636363FE");
        foo := test(x"0000000000000000000000000000000D");
        wait for delay;
        foo := as(x"636363636363636363636363636363D7");
        foo := test(x"0000000000000000000000000000000E");
        wait for delay;
        foo := as(x"636363636363636363636363636363AB");
        foo := test(x"0000000000000000000000000000000F");
        wait for delay;
        foo := as(x"63636363636363636363636363636376");
        foo := test(x"00000000000000000000000000000010");
        wait for delay;
        foo := as(x"636363636363636363636363636363CA");
        foo := test(x"00000000000000000000000000000011");
        wait for delay;
        foo := as(x"63636363636363636363636363636382");
        foo := test(x"00000000000000000000000000000012");
        wait for delay;
        foo := as(x"636363636363636363636363636363C9");
        foo := test(x"00000000000000000000000000000013");
        wait for delay;
        foo := as(x"6363636363636363636363636363637D");
        foo := test(x"00000000000000000000000000000014");
        wait for delay;
        foo := as(x"636363636363636363636363636363FA");
        foo := test(x"00000000000000000000000000000015");
        wait for delay;
        foo := as(x"63636363636363636363636363636359");
        foo := test(x"00000000000000000000000000000016");
        wait for delay;
        foo := as(x"63636363636363636363636363636347");
        foo := test(x"00000000000000000000000000000017");
        wait for delay;
        foo := as(x"636363636363636363636363636363F0");
        foo := test(x"00000000000000000000000000000018");
        wait for delay;
        foo := as(x"636363636363636363636363636363AD");
        foo := test(x"00000000000000000000000000000019");
        wait for delay;
        foo := as(x"636363636363636363636363636363D4");
        foo := test(x"0000000000000000000000000000001A");
        wait for delay;
        foo := as(x"636363636363636363636363636363A2");
        foo := test(x"0000000000000000000000000000001B");
        wait for delay;
        foo := as(x"636363636363636363636363636363AF");
        foo := test(x"0000000000000000000000000000001C");
        wait for delay;
        foo := as(x"6363636363636363636363636363639C");
        foo := test(x"0000000000000000000000000000001D");
        wait for delay;
        foo := as(x"636363636363636363636363636363A4");
        foo := test(x"0000000000000000000000000000001E");
        wait for delay;
        foo := as(x"63636363636363636363636363636372");
        foo := test(x"0000000000000000000000000000001F");
        wait for delay;
        foo := as(x"636363636363636363636363636363C0");
        foo := test(x"00000000000000000000000000000020");
        wait for delay;
        foo := as(x"636363636363636363636363636363B7");
        foo := test(x"00000000000000000000000000000021");
        wait for delay;
        foo := as(x"636363636363636363636363636363FD");
        foo := test(x"00000000000000000000000000000022");
        wait for delay;
        foo := as(x"63636363636363636363636363636393");
        foo := test(x"00000000000000000000000000000023");
        wait for delay;
        foo := as(x"63636363636363636363636363636326");
        foo := test(x"00000000000000000000000000000024");
        wait for delay;
        foo := as(x"63636363636363636363636363636336");
        foo := test(x"00000000000000000000000000000025");
        wait for delay;
        foo := as(x"6363636363636363636363636363633F");
        foo := test(x"00000000000000000000000000000026");
        wait for delay;
        foo := as(x"636363636363636363636363636363F7");
        foo := test(x"00000000000000000000000000000027");
        wait for delay;
        foo := as(x"636363636363636363636363636363CC");
        foo := test(x"00000000000000000000000000000028");
        wait for delay;
        foo := as(x"63636363636363636363636363636334");
        foo := test(x"00000000000000000000000000000029");
        wait for delay;
        foo := as(x"636363636363636363636363636363A5");
        foo := test(x"0000000000000000000000000000002A");
        wait for delay;
        foo := as(x"636363636363636363636363636363E5");
        foo := test(x"0000000000000000000000000000002B");
        wait for delay;
        foo := as(x"636363636363636363636363636363F1");
        foo := test(x"0000000000000000000000000000002C");
        wait for delay;
        foo := as(x"63636363636363636363636363636371");
        foo := test(x"0000000000000000000000000000002D");
        wait for delay;
        foo := as(x"636363636363636363636363636363D8");
        foo := test(x"0000000000000000000000000000002E");
        wait for delay;
        foo := as(x"63636363636363636363636363636331");
        foo := test(x"0000000000000000000000000000002F");
        wait for delay;
        foo := as(x"63636363636363636363636363636315");
        foo := test(x"00000000000000000000000000000030");
        wait for delay;
        foo := as(x"63636363636363636363636363636304");
        foo := test(x"00000000000000000000000000000031");
        wait for delay;
        foo := as(x"636363636363636363636363636363C7");
        foo := test(x"00000000000000000000000000000032");
        wait for delay;
        foo := as(x"63636363636363636363636363636323");
        foo := test(x"00000000000000000000000000000033");
        wait for delay;
        foo := as(x"636363636363636363636363636363C3");
        foo := test(x"00000000000000000000000000000034");
        wait for delay;
        foo := as(x"63636363636363636363636363636318");
        foo := test(x"00000000000000000000000000000035");
        wait for delay;
        foo := as(x"63636363636363636363636363636396");
        foo := test(x"00000000000000000000000000000036");
        wait for delay;
        foo := as(x"63636363636363636363636363636305");
        foo := test(x"00000000000000000000000000000037");
        wait for delay;
        foo := as(x"6363636363636363636363636363639A");
        foo := test(x"00000000000000000000000000000038");
        wait for delay;
        foo := as(x"63636363636363636363636363636307");
        foo := test(x"00000000000000000000000000000039");
        wait for delay;
        foo := as(x"63636363636363636363636363636312");
        foo := test(x"0000000000000000000000000000003A");
        wait for delay;
        foo := as(x"63636363636363636363636363636380");
        foo := test(x"0000000000000000000000000000003B");
        wait for delay;
        foo := as(x"636363636363636363636363636363E2");
        foo := test(x"0000000000000000000000000000003C");
        wait for delay;
        foo := as(x"636363636363636363636363636363EB");
        foo := test(x"0000000000000000000000000000003D");
        wait for delay;
        foo := as(x"63636363636363636363636363636327");
        foo := test(x"0000000000000000000000000000003E");
        wait for delay;
        foo := as(x"636363636363636363636363636363B2");
        foo := test(x"0000000000000000000000000000003F");
        wait for delay;
        foo := as(x"63636363636363636363636363636375");
        foo := test(x"00000000000000000000000000000040");
        wait for delay;
        foo := as(x"63636363636363636363636363636309");
        foo := test(x"00000000000000000000000000000041");
        wait for delay;
        foo := as(x"63636363636363636363636363636383");
        foo := test(x"00000000000000000000000000000042");
        wait for delay;
        foo := as(x"6363636363636363636363636363632C");
        foo := test(x"00000000000000000000000000000043");
        wait for delay;
        foo := as(x"6363636363636363636363636363631A");
        foo := test(x"00000000000000000000000000000044");
        wait for delay;
        foo := as(x"6363636363636363636363636363631B");
        foo := test(x"00000000000000000000000000000045");
        wait for delay;
        foo := as(x"6363636363636363636363636363636E");
        foo := test(x"00000000000000000000000000000046");
        wait for delay;
        foo := as(x"6363636363636363636363636363635A");
        foo := test(x"00000000000000000000000000000047");
        wait for delay;
        foo := as(x"636363636363636363636363636363A0");
        foo := test(x"00000000000000000000000000000048");
        wait for delay;
        foo := as(x"63636363636363636363636363636352");
        foo := test(x"00000000000000000000000000000049");
        wait for delay;
        foo := as(x"6363636363636363636363636363633B");
        foo := test(x"0000000000000000000000000000004A");
        wait for delay;
        foo := as(x"636363636363636363636363636363D6");
        foo := test(x"0000000000000000000000000000004B");
        wait for delay;
        foo := as(x"636363636363636363636363636363B3");
        foo := test(x"0000000000000000000000000000004C");
        wait for delay;
        foo := as(x"63636363636363636363636363636329");
        foo := test(x"0000000000000000000000000000004D");
        wait for delay;
        foo := as(x"636363636363636363636363636363E3");
        foo := test(x"0000000000000000000000000000004E");
        wait for delay;
        foo := as(x"6363636363636363636363636363632F");
        foo := test(x"0000000000000000000000000000004F");
        wait for delay;
        foo := as(x"63636363636363636363636363636384");
        foo := test(x"00000000000000000000000000000050");
        wait for delay;
        foo := as(x"63636363636363636363636363636353");
        foo := test(x"00000000000000000000000000000051");
        wait for delay;
        foo := as(x"636363636363636363636363636363D1");
        foo := test(x"00000000000000000000000000000052");
        wait for delay;
        foo := as(x"63636363636363636363636363636300");
        foo := test(x"00000000000000000000000000000053");
        wait for delay;
        foo := as(x"636363636363636363636363636363ED");
        foo := test(x"00000000000000000000000000000054");
        wait for delay;
        foo := as(x"63636363636363636363636363636320");
        foo := test(x"00000000000000000000000000000055");
        wait for delay;
        foo := as(x"636363636363636363636363636363FC");
        foo := test(x"00000000000000000000000000000056");
        wait for delay;
        foo := as(x"636363636363636363636363636363B1");
        foo := test(x"00000000000000000000000000000057");
        wait for delay;
        foo := as(x"6363636363636363636363636363635B");
        foo := test(x"00000000000000000000000000000058");
        wait for delay;
        foo := as(x"6363636363636363636363636363636A");
        foo := test(x"00000000000000000000000000000059");
        wait for delay;
        foo := as(x"636363636363636363636363636363CB");
        foo := test(x"0000000000000000000000000000005A");
        wait for delay;
        foo := as(x"636363636363636363636363636363BE");
        foo := test(x"0000000000000000000000000000005B");
        wait for delay;
        foo := as(x"63636363636363636363636363636339");
        foo := test(x"0000000000000000000000000000005C");
        wait for delay;
        foo := as(x"6363636363636363636363636363634A");
        foo := test(x"0000000000000000000000000000005D");
        wait for delay;
        foo := as(x"6363636363636363636363636363634C");
        foo := test(x"0000000000000000000000000000005E");
        wait for delay;
        foo := as(x"63636363636363636363636363636358");
        foo := test(x"0000000000000000000000000000005F");
        wait for delay;
        foo := as(x"636363636363636363636363636363CF");
        foo := test(x"00000000000000000000000000000060");
        wait for delay;
        foo := as(x"636363636363636363636363636363D0");
        foo := test(x"00000000000000000000000000000061");
        wait for delay;
        foo := as(x"636363636363636363636363636363EF");
        foo := test(x"00000000000000000000000000000062");
        wait for delay;
        foo := as(x"636363636363636363636363636363AA");
        foo := test(x"00000000000000000000000000000063");
        wait for delay;
        foo := as(x"636363636363636363636363636363FB");
        foo := test(x"00000000000000000000000000000064");
        wait for delay;
        foo := as(x"63636363636363636363636363636343");
        foo := test(x"00000000000000000000000000000065");
        wait for delay;
        foo := as(x"6363636363636363636363636363634D");
        foo := test(x"00000000000000000000000000000066");
        wait for delay;
        foo := as(x"63636363636363636363636363636333");
        foo := test(x"00000000000000000000000000000067");
        wait for delay;
        foo := as(x"63636363636363636363636363636385");
        foo := test(x"00000000000000000000000000000068");
        wait for delay;
        foo := as(x"63636363636363636363636363636345");
        foo := test(x"00000000000000000000000000000069");
        wait for delay;
        foo := as(x"636363636363636363636363636363F9");
        foo := test(x"0000000000000000000000000000006A");
        wait for delay;
        foo := as(x"63636363636363636363636363636302");
        foo := test(x"0000000000000000000000000000006B");
        wait for delay;
        foo := as(x"6363636363636363636363636363637F");
        foo := test(x"0000000000000000000000000000006C");
        wait for delay;
        foo := as(x"63636363636363636363636363636350");
        foo := test(x"0000000000000000000000000000006D");
        wait for delay;
        foo := as(x"6363636363636363636363636363633C");
        foo := test(x"0000000000000000000000000000006E");
        wait for delay;
        foo := as(x"6363636363636363636363636363639F");
        foo := test(x"0000000000000000000000000000006F");
        wait for delay;
        foo := as(x"636363636363636363636363636363A8");
        foo := test(x"00000000000000000000000000000070");
        wait for delay;
        foo := as(x"63636363636363636363636363636351");
        foo := test(x"00000000000000000000000000000071");
        wait for delay;
        foo := as(x"636363636363636363636363636363A3");
        foo := test(x"00000000000000000000000000000072");
        wait for delay;
        foo := as(x"63636363636363636363636363636340");
        foo := test(x"00000000000000000000000000000073");
        wait for delay;
        foo := as(x"6363636363636363636363636363638F");
        foo := test(x"00000000000000000000000000000074");
        wait for delay;
        foo := as(x"63636363636363636363636363636392");
        foo := test(x"00000000000000000000000000000075");
        wait for delay;
        foo := as(x"6363636363636363636363636363639D");
        foo := test(x"00000000000000000000000000000076");
        wait for delay;
        foo := as(x"63636363636363636363636363636338");
        foo := test(x"00000000000000000000000000000077");
        wait for delay;
        foo := as(x"636363636363636363636363636363F5");
        foo := test(x"00000000000000000000000000000078");
        wait for delay;
        foo := as(x"636363636363636363636363636363BC");
        foo := test(x"00000000000000000000000000000079");
        wait for delay;
        foo := as(x"636363636363636363636363636363B6");
        foo := test(x"0000000000000000000000000000007A");
        wait for delay;
        foo := as(x"636363636363636363636363636363DA");
        foo := test(x"0000000000000000000000000000007B");
        wait for delay;
        foo := as(x"63636363636363636363636363636321");
        foo := test(x"0000000000000000000000000000007C");
        wait for delay;
        foo := as(x"63636363636363636363636363636310");
        foo := test(x"0000000000000000000000000000007D");
        wait for delay;
        foo := as(x"636363636363636363636363636363FF");
        foo := test(x"0000000000000000000000000000007E");
        wait for delay;
        foo := as(x"636363636363636363636363636363F3");
        foo := test(x"0000000000000000000000000000007F");
        wait for delay;
        foo := as(x"636363636363636363636363636363D2");
        foo := test(x"00000000000000000000000000000080");
        wait for delay;
        foo := as(x"636363636363636363636363636363CD");
        foo := test(x"00000000000000000000000000000081");
        wait for delay;
        foo := as(x"6363636363636363636363636363630C");
        foo := test(x"00000000000000000000000000000082");
        wait for delay;
        foo := as(x"63636363636363636363636363636313");
        foo := test(x"00000000000000000000000000000083");
        wait for delay;
        foo := as(x"636363636363636363636363636363EC");
        foo := test(x"00000000000000000000000000000084");
        wait for delay;
        foo := as(x"6363636363636363636363636363635F");
        foo := test(x"00000000000000000000000000000085");
        wait for delay;
        foo := as(x"63636363636363636363636363636397");
        foo := test(x"00000000000000000000000000000086");
        wait for delay;
        foo := as(x"63636363636363636363636363636344");
        foo := test(x"00000000000000000000000000000087");
        wait for delay;
        foo := as(x"63636363636363636363636363636317");
        foo := test(x"00000000000000000000000000000088");
        wait for delay;
        foo := as(x"636363636363636363636363636363C4");
        foo := test(x"00000000000000000000000000000089");
        wait for delay;
        foo := as(x"636363636363636363636363636363A7");
        foo := test(x"0000000000000000000000000000008A");
        wait for delay;
        foo := as(x"6363636363636363636363636363637E");
        foo := test(x"0000000000000000000000000000008B");
        wait for delay;
        foo := as(x"6363636363636363636363636363633D");
        foo := test(x"0000000000000000000000000000008C");
        wait for delay;
        foo := as(x"63636363636363636363636363636364");
        foo := test(x"0000000000000000000000000000008D");
        wait for delay;
        foo := as(x"6363636363636363636363636363635D");
        foo := test(x"0000000000000000000000000000008E");
        wait for delay;
        foo := as(x"63636363636363636363636363636319");
        foo := test(x"0000000000000000000000000000008F");
        wait for delay;
        foo := as(x"63636363636363636363636363636373");
        foo := test(x"00000000000000000000000000000090");
        wait for delay;
        foo := as(x"63636363636363636363636363636360");
        foo := test(x"00000000000000000000000000000091");
        wait for delay;
        foo := as(x"63636363636363636363636363636381");
        foo := test(x"00000000000000000000000000000092");
        wait for delay;
        foo := as(x"6363636363636363636363636363634F");
        foo := test(x"00000000000000000000000000000093");
        wait for delay;
        foo := as(x"636363636363636363636363636363DC");
        foo := test(x"00000000000000000000000000000094");
        wait for delay;
        foo := as(x"63636363636363636363636363636322");
        foo := test(x"00000000000000000000000000000095");
        wait for delay;
        foo := as(x"6363636363636363636363636363632A");
        foo := test(x"00000000000000000000000000000096");
        wait for delay;
        foo := as(x"63636363636363636363636363636390");
        foo := test(x"00000000000000000000000000000097");
        wait for delay;
        foo := as(x"63636363636363636363636363636388");
        foo := test(x"00000000000000000000000000000098");
        wait for delay;
        foo := as(x"63636363636363636363636363636346");
        foo := test(x"00000000000000000000000000000099");
        wait for delay;
        foo := as(x"636363636363636363636363636363EE");
        foo := test(x"0000000000000000000000000000009A");
        wait for delay;
        foo := as(x"636363636363636363636363636363B8");
        foo := test(x"0000000000000000000000000000009B");
        wait for delay;
        foo := as(x"63636363636363636363636363636314");
        foo := test(x"0000000000000000000000000000009C");
        wait for delay;
        foo := as(x"636363636363636363636363636363DE");
        foo := test(x"0000000000000000000000000000009D");
        wait for delay;
        foo := as(x"6363636363636363636363636363635E");
        foo := test(x"0000000000000000000000000000009E");
        wait for delay;
        foo := as(x"6363636363636363636363636363630B");
        foo := test(x"0000000000000000000000000000009F");
        wait for delay;
        foo := as(x"636363636363636363636363636363DB");
        foo := test(x"000000000000000000000000000000A0");
        wait for delay;
        foo := as(x"636363636363636363636363636363E0");
        foo := test(x"000000000000000000000000000000A1");
        wait for delay;
        foo := as(x"63636363636363636363636363636332");
        foo := test(x"000000000000000000000000000000A2");
        wait for delay;
        foo := as(x"6363636363636363636363636363633A");
        foo := test(x"000000000000000000000000000000A3");
        wait for delay;
        foo := as(x"6363636363636363636363636363630A");
        foo := test(x"000000000000000000000000000000A4");
        wait for delay;
        foo := as(x"63636363636363636363636363636349");
        foo := test(x"000000000000000000000000000000A5");
        wait for delay;
        foo := as(x"63636363636363636363636363636306");
        foo := test(x"000000000000000000000000000000A6");
        wait for delay;
        foo := as(x"63636363636363636363636363636324");
        foo := test(x"000000000000000000000000000000A7");
        wait for delay;
        foo := as(x"6363636363636363636363636363635C");
        foo := test(x"000000000000000000000000000000A8");
        wait for delay;
        foo := as(x"636363636363636363636363636363C2");
        foo := test(x"000000000000000000000000000000A9");
        wait for delay;
        foo := as(x"636363636363636363636363636363D3");
        foo := test(x"000000000000000000000000000000AA");
        wait for delay;
        foo := as(x"636363636363636363636363636363AC");
        foo := test(x"000000000000000000000000000000AB");
        wait for delay;
        foo := as(x"63636363636363636363636363636362");
        foo := test(x"000000000000000000000000000000AC");
        wait for delay;
        foo := as(x"63636363636363636363636363636391");
        foo := test(x"000000000000000000000000000000AD");
        wait for delay;
        foo := as(x"63636363636363636363636363636395");
        foo := test(x"000000000000000000000000000000AE");
        wait for delay;
        foo := as(x"636363636363636363636363636363E4");
        foo := test(x"000000000000000000000000000000AF");
        wait for delay;
        foo := as(x"63636363636363636363636363636379");
        foo := test(x"000000000000000000000000000000B0");
        wait for delay;
        foo := as(x"636363636363636363636363636363E7");
        foo := test(x"000000000000000000000000000000B1");
        wait for delay;
        foo := as(x"636363636363636363636363636363C8");
        foo := test(x"000000000000000000000000000000B2");
        wait for delay;
        foo := as(x"63636363636363636363636363636337");
        foo := test(x"000000000000000000000000000000B3");
        wait for delay;
        foo := as(x"6363636363636363636363636363636D");
        foo := test(x"000000000000000000000000000000B4");
        wait for delay;
        foo := as(x"6363636363636363636363636363638D");
        foo := test(x"000000000000000000000000000000B5");
        wait for delay;
        foo := as(x"636363636363636363636363636363D5");
        foo := test(x"000000000000000000000000000000B6");
        wait for delay;
        foo := as(x"6363636363636363636363636363634E");
        foo := test(x"000000000000000000000000000000B7");
        wait for delay;
        foo := as(x"636363636363636363636363636363A9");
        foo := test(x"000000000000000000000000000000B8");
        wait for delay;
        foo := as(x"6363636363636363636363636363636C");
        foo := test(x"000000000000000000000000000000B9");
        wait for delay;
        foo := as(x"63636363636363636363636363636356");
        foo := test(x"000000000000000000000000000000BA");
        wait for delay;
        foo := as(x"636363636363636363636363636363F4");
        foo := test(x"000000000000000000000000000000BB");
        wait for delay;
        foo := as(x"636363636363636363636363636363EA");
        foo := test(x"000000000000000000000000000000BC");
        wait for delay;
        foo := as(x"63636363636363636363636363636365");
        foo := test(x"000000000000000000000000000000BD");
        wait for delay;
        foo := as(x"6363636363636363636363636363637A");
        foo := test(x"000000000000000000000000000000BE");
        wait for delay;
        foo := as(x"636363636363636363636363636363AE");
        foo := test(x"000000000000000000000000000000BF");
        wait for delay;
        foo := as(x"63636363636363636363636363636308");
        foo := test(x"000000000000000000000000000000C0");
        wait for delay;
        foo := as(x"636363636363636363636363636363BA");
        foo := test(x"000000000000000000000000000000C1");
        wait for delay;
        foo := as(x"63636363636363636363636363636378");
        foo := test(x"000000000000000000000000000000C2");
        wait for delay;
        foo := as(x"63636363636363636363636363636325");
        foo := test(x"000000000000000000000000000000C3");
        wait for delay;
        foo := as(x"6363636363636363636363636363632E");
        foo := test(x"000000000000000000000000000000C4");
        wait for delay;
        foo := as(x"6363636363636363636363636363631C");
        foo := test(x"000000000000000000000000000000C5");
        wait for delay;
        foo := as(x"636363636363636363636363636363A6");
        foo := test(x"000000000000000000000000000000C6");
        wait for delay;
        foo := as(x"636363636363636363636363636363B4");
        foo := test(x"000000000000000000000000000000C7");
        wait for delay;
        foo := as(x"636363636363636363636363636363C6");
        foo := test(x"000000000000000000000000000000C8");
        wait for delay;
        foo := as(x"636363636363636363636363636363E8");
        foo := test(x"000000000000000000000000000000C9");
        wait for delay;
        foo := as(x"636363636363636363636363636363DD");
        foo := test(x"000000000000000000000000000000CA");
        wait for delay;
        foo := as(x"63636363636363636363636363636374");
        foo := test(x"000000000000000000000000000000CB");
        wait for delay;
        foo := as(x"6363636363636363636363636363631F");
        foo := test(x"000000000000000000000000000000CC");
        wait for delay;
        foo := as(x"6363636363636363636363636363634B");
        foo := test(x"000000000000000000000000000000CD");
        wait for delay;
        foo := as(x"636363636363636363636363636363BD");
        foo := test(x"000000000000000000000000000000CE");
        wait for delay;
        foo := as(x"6363636363636363636363636363638B");
        foo := test(x"000000000000000000000000000000CF");
        wait for delay;
        foo := as(x"6363636363636363636363636363638A");
        foo := test(x"000000000000000000000000000000D0");
        wait for delay;
        foo := as(x"63636363636363636363636363636370");
        foo := test(x"000000000000000000000000000000D1");
        wait for delay;
        foo := as(x"6363636363636363636363636363633E");
        foo := test(x"000000000000000000000000000000D2");
        wait for delay;
        foo := as(x"636363636363636363636363636363B5");
        foo := test(x"000000000000000000000000000000D3");
        wait for delay;
        foo := as(x"63636363636363636363636363636366");
        foo := test(x"000000000000000000000000000000D4");
        wait for delay;
        foo := as(x"63636363636363636363636363636348");
        foo := test(x"000000000000000000000000000000D5");
        wait for delay;
        foo := as(x"63636363636363636363636363636303");
        foo := test(x"000000000000000000000000000000D6");
        wait for delay;
        foo := as(x"636363636363636363636363636363F6");
        foo := test(x"000000000000000000000000000000D7");
        wait for delay;
        foo := as(x"6363636363636363636363636363630E");
        foo := test(x"000000000000000000000000000000D8");
        wait for delay;
        foo := as(x"63636363636363636363636363636361");
        foo := test(x"000000000000000000000000000000D9");
        wait for delay;
        foo := as(x"63636363636363636363636363636335");
        foo := test(x"000000000000000000000000000000DA");
        wait for delay;
        foo := as(x"63636363636363636363636363636357");
        foo := test(x"000000000000000000000000000000DB");
        wait for delay;
        foo := as(x"636363636363636363636363636363B9");
        foo := test(x"000000000000000000000000000000DC");
        wait for delay;
        foo := as(x"63636363636363636363636363636386");
        foo := test(x"000000000000000000000000000000DD");
        wait for delay;
        foo := as(x"636363636363636363636363636363C1");
        foo := test(x"000000000000000000000000000000DE");
        wait for delay;
        foo := as(x"6363636363636363636363636363631D");
        foo := test(x"000000000000000000000000000000DF");
        wait for delay;
        foo := as(x"6363636363636363636363636363639E");
        foo := test(x"000000000000000000000000000000E0");
        wait for delay;
        foo := as(x"636363636363636363636363636363E1");
        foo := test(x"000000000000000000000000000000E1");
        wait for delay;
        foo := as(x"636363636363636363636363636363F8");
        foo := test(x"000000000000000000000000000000E2");
        wait for delay;
        foo := as(x"63636363636363636363636363636398");
        foo := test(x"000000000000000000000000000000E3");
        wait for delay;
        foo := as(x"63636363636363636363636363636311");
        foo := test(x"000000000000000000000000000000E4");
        wait for delay;
        foo := as(x"63636363636363636363636363636369");
        foo := test(x"000000000000000000000000000000E5");
        wait for delay;
        foo := as(x"636363636363636363636363636363D9");
        foo := test(x"000000000000000000000000000000E6");
        wait for delay;
        foo := as(x"6363636363636363636363636363638E");
        foo := test(x"000000000000000000000000000000E7");
        wait for delay;
        foo := as(x"63636363636363636363636363636394");
        foo := test(x"000000000000000000000000000000E8");
        wait for delay;
        foo := as(x"6363636363636363636363636363639B");
        foo := test(x"000000000000000000000000000000E9");
        wait for delay;
        foo := as(x"6363636363636363636363636363631E");
        foo := test(x"000000000000000000000000000000EA");
        wait for delay;
        foo := as(x"63636363636363636363636363636387");
        foo := test(x"000000000000000000000000000000EB");
        wait for delay;
        foo := as(x"636363636363636363636363636363E9");
        foo := test(x"000000000000000000000000000000EC");
        wait for delay;
        foo := as(x"636363636363636363636363636363CE");
        foo := test(x"000000000000000000000000000000ED");
        wait for delay;
        foo := as(x"63636363636363636363636363636355");
        foo := test(x"000000000000000000000000000000EE");
        wait for delay;
        foo := as(x"63636363636363636363636363636328");
        foo := test(x"000000000000000000000000000000EF");
        wait for delay;
        foo := as(x"636363636363636363636363636363DF");
        foo := test(x"000000000000000000000000000000F0");
        wait for delay;
        foo := as(x"6363636363636363636363636363638C");
        foo := test(x"000000000000000000000000000000F1");
        wait for delay;
        foo := as(x"636363636363636363636363636363A1");
        foo := test(x"000000000000000000000000000000F2");
        wait for delay;
        foo := as(x"63636363636363636363636363636389");
        foo := test(x"000000000000000000000000000000F3");
        wait for delay;
        foo := as(x"6363636363636363636363636363630D");
        foo := test(x"000000000000000000000000000000F4");
        wait for delay;
        foo := as(x"636363636363636363636363636363BF");
        foo := test(x"000000000000000000000000000000F5");
        wait for delay;
        foo := as(x"636363636363636363636363636363E6");
        foo := test(x"000000000000000000000000000000F6");
        wait for delay;
        foo := as(x"63636363636363636363636363636342");
        foo := test(x"000000000000000000000000000000F7");
        wait for delay;
        foo := as(x"63636363636363636363636363636368");
        foo := test(x"000000000000000000000000000000F8");
        wait for delay;
        foo := as(x"63636363636363636363636363636341");
        foo := test(x"000000000000000000000000000000F9");
        wait for delay;
        foo := as(x"63636363636363636363636363636399");
        foo := test(x"000000000000000000000000000000FA");
        wait for delay;
        foo := as(x"6363636363636363636363636363632D");
        foo := test(x"000000000000000000000000000000FB");
        wait for delay;
        foo := as(x"6363636363636363636363636363630F");
        foo := test(x"000000000000000000000000000000FC");
        wait for delay;
        foo := as(x"636363636363636363636363636363B0");
        foo := test(x"000000000000000000000000000000FD");
        wait for delay;
        foo := as(x"63636363636363636363636363636354");
        foo := test(x"000000000000000000000000000000FE");
        wait for delay;
        foo := as(x"636363636363636363636363636363BB");
        foo := test(x"000000000000000000000000000000FF");
        wait for delay;
        foo := as(x"63636363636363636363636363636316");
        
    end process;
end tb;
