LIBRARY ieee;
USE ieee.std_logic_1164.all;

entity InverseSBoxTb is
end InverseSBoxTb;

architecture ISBoxTb of InverseSBoxTb is
  component InverseSubstituteBox
    port
    (
      data_in : in std_logic_vector(127 downto 0);
      data_out : out std_logic_Vector(127 downto 0)
    );
  end component;

  signal data_in  : std_logic_vector(127 downto 0);
  signal data_out : std_logic_Vector(127 downto 0);

  signal delay : time := 20 ns;

  begin
    InverseSBoxPort : InverseSubstituteBox port map (
      data_in => data_in,
      data_out => data_out
    );

    process
    begin
      data_in <= x"00000000000000000000000000000000";
      wait for delay;
      assert data_out = x"52525252525252525252525252525252" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000001";
      wait for delay;
      assert data_out = x"52525252525252525252525252525209" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000002";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526A" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000003";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D5" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000004";
      wait for delay;
      assert data_out = x"52525252525252525252525252525230" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000005";
      wait for delay;
      assert data_out = x"52525252525252525252525252525236" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000006";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A5" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000007";
      wait for delay;
      assert data_out = x"52525252525252525252525252525238" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000008";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BF" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000009";
      wait for delay;
      assert data_out = x"52525252525252525252525252525240" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000A";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A3" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000B";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529E" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000C";
      wait for delay;
      assert data_out = x"52525252525252525252525252525281" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000D";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F3" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D7" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000000F";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FB" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000010";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527C" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000011";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E3" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000012";
      wait for delay;
      assert data_out = x"52525252525252525252525252525239" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000013";
      wait for delay;
      assert data_out = x"52525252525252525252525252525282" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000014";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529B" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000015";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522F" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000016";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FF" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000017";
      wait for delay;
      assert data_out = x"52525252525252525252525252525287" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000018";
      wait for delay;
      assert data_out = x"52525252525252525252525252525234" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000019";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528E" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001A";
      wait for delay;
      assert data_out = x"52525252525252525252525252525243" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001B";
      wait for delay;
      assert data_out = x"52525252525252525252525252525244" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001C";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C4" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001D";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DE" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E9" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000001F";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CB" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000020";
      wait for delay;
      assert data_out = x"52525252525252525252525252525254" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000021";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527B" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000022";
      wait for delay;
      assert data_out = x"52525252525252525252525252525294" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000023";
      wait for delay;
      assert data_out = x"52525252525252525252525252525232" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000024";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A6" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000025";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C2" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000026";
      wait for delay;
      assert data_out = x"52525252525252525252525252525223" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000027";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523D" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000028";
      wait for delay;
      assert data_out = x"525252525252525252525252525252EE" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000029";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524C" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002A";
      wait for delay;
      assert data_out = x"52525252525252525252525252525295" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002B";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520B" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002C";
      wait for delay;
      assert data_out = x"52525252525252525252525252525242" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002D";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FA" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C3" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000002F";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524E" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000030";
      wait for delay;
      assert data_out = x"52525252525252525252525252525208" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000031";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522E" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000032";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A1" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000033";
      wait for delay;
      assert data_out = x"52525252525252525252525252525266" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000034";
      wait for delay;
      assert data_out = x"52525252525252525252525252525228" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000035";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D9" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000036";
      wait for delay;
      assert data_out = x"52525252525252525252525252525224" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000037";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B2" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000038";
      wait for delay;
      assert data_out = x"52525252525252525252525252525276" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000039";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525B" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003A";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A2" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003B";
      wait for delay;
      assert data_out = x"52525252525252525252525252525249" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003C";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526D" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003D";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528B" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D1" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000003F";
      wait for delay;
      assert data_out = x"52525252525252525252525252525225" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000040";
      wait for delay;
      assert data_out = x"52525252525252525252525252525272" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000041";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F8" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000042";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F6" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000043";
      wait for delay;
      assert data_out = x"52525252525252525252525252525264" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000044";
      wait for delay;
      assert data_out = x"52525252525252525252525252525286" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000045";
      wait for delay;
      assert data_out = x"52525252525252525252525252525268" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000046";
      wait for delay;
      assert data_out = x"52525252525252525252525252525298" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000047";
      wait for delay;
      assert data_out = x"52525252525252525252525252525216" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000048";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D4" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000049";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A4" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004A";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525C" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004B";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CC" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004C";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525D" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004D";
      wait for delay;
      assert data_out = x"52525252525252525252525252525265" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B6" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000004F";
      wait for delay;
      assert data_out = x"52525252525252525252525252525292" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000050";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526C" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000051";
      wait for delay;
      assert data_out = x"52525252525252525252525252525270" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000052";
      wait for delay;
      assert data_out = x"52525252525252525252525252525248" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000053";
      wait for delay;
      assert data_out = x"52525252525252525252525252525250" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000054";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FD" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000055";
      wait for delay;
      assert data_out = x"525252525252525252525252525252ED" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000056";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B9" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000057";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DA" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000058";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525E" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000059";
      wait for delay;
      assert data_out = x"52525252525252525252525252525215" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005A";
      wait for delay;
      assert data_out = x"52525252525252525252525252525246" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005B";
      wait for delay;
      assert data_out = x"52525252525252525252525252525257" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005C";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A7" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005D";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528D" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005E";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529D" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000005F";
      wait for delay;
      assert data_out = x"52525252525252525252525252525284" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000060";
      wait for delay;
      assert data_out = x"52525252525252525252525252525290" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000061";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D8" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000062";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AB" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000063";
      wait for delay;
      assert data_out = x"52525252525252525252525252525200" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000064";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528C" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000065";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BC" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000066";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D3" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000067";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520A" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000068";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F7" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000069";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E4" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006A";
      wait for delay;
      assert data_out = x"52525252525252525252525252525258" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006B";
      wait for delay;
      assert data_out = x"52525252525252525252525252525205" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006C";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B8" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006D";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B3" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006E";
      wait for delay;
      assert data_out = x"52525252525252525252525252525245" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000006F";
      wait for delay;
      assert data_out = x"52525252525252525252525252525206" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000070";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D0" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000071";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522C" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000072";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521E" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000073";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528F" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000074";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CA" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000075";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523F" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000076";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520F" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000077";
      wait for delay;
      assert data_out = x"52525252525252525252525252525202" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000078";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C1" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000079";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AF" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007A";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BD" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007B";
      wait for delay;
      assert data_out = x"52525252525252525252525252525203" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007C";
      wait for delay;
      assert data_out = x"52525252525252525252525252525201" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007D";
      wait for delay;
      assert data_out = x"52525252525252525252525252525213" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007E";
      wait for delay;
      assert data_out = x"5252525252525252525252525252528A" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000007F";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526B" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000080";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523A" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000081";
      wait for delay;
      assert data_out = x"52525252525252525252525252525291" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000082";
      wait for delay;
      assert data_out = x"52525252525252525252525252525211" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000083";
      wait for delay;
      assert data_out = x"52525252525252525252525252525241" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000084";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524F" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000085";
      wait for delay;
      assert data_out = x"52525252525252525252525252525267" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000086";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DC" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000087";
      wait for delay;
      assert data_out = x"525252525252525252525252525252EA" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000088";
      wait for delay;
      assert data_out = x"52525252525252525252525252525297" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000089";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F2" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008A";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CF" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008B";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CE" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008C";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F0" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008D";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B4" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E6" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000008F";
      wait for delay;
      assert data_out = x"52525252525252525252525252525273" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000090";
      wait for delay;
      assert data_out = x"52525252525252525252525252525296" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000091";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AC" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000092";
      wait for delay;
      assert data_out = x"52525252525252525252525252525274" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000093";
      wait for delay;
      assert data_out = x"52525252525252525252525252525222" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000094";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E7" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000095";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AD" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000096";
      wait for delay;
      assert data_out = x"52525252525252525252525252525235" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000097";
      wait for delay;
      assert data_out = x"52525252525252525252525252525285" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000098";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E2" report "Inverse SBox wrong" severity error;
      data_in <= x"00000000000000000000000000000099";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F9" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009A";
      wait for delay;
      assert data_out = x"52525252525252525252525252525237" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009B";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E8" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009C";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521C" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009D";
      wait for delay;
      assert data_out = x"52525252525252525252525252525275" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009E";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DF" report "Inverse SBox wrong" severity error;
      data_in <= x"0000000000000000000000000000009F";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526E" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A0";
      wait for delay;
      assert data_out = x"52525252525252525252525252525247" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A1";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F1" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A2";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A3";
      wait for delay;
      assert data_out = x"52525252525252525252525252525271" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A4";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521D" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A5";
      wait for delay;
      assert data_out = x"52525252525252525252525252525229" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A6";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C5" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A7";
      wait for delay;
      assert data_out = x"52525252525252525252525252525289" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A8";
      wait for delay;
      assert data_out = x"5252525252525252525252525252526F" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000A9";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B7" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AA";
      wait for delay;
      assert data_out = x"52525252525252525252525252525262" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AB";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520E" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AC";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AA" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AD";
      wait for delay;
      assert data_out = x"52525252525252525252525252525218" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AE";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BE" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000AF";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521B" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B0";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FC" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B1";
      wait for delay;
      assert data_out = x"52525252525252525252525252525256" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B2";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523E" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B3";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524B" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B4";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C6" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B5";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D2" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B6";
      wait for delay;
      assert data_out = x"52525252525252525252525252525279" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B7";
      wait for delay;
      assert data_out = x"52525252525252525252525252525220" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B8";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000B9";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DB" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BA";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C0" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BB";
      wait for delay;
      assert data_out = x"525252525252525252525252525252FE" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BC";
      wait for delay;
      assert data_out = x"52525252525252525252525252525278" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BD";
      wait for delay;
      assert data_out = x"525252525252525252525252525252CD" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BE";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000BF";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F4" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C0";
      wait for delay;
      assert data_out = x"5252525252525252525252525252521F" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C1";
      wait for delay;
      assert data_out = x"525252525252525252525252525252DD" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C2";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A8" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C3";
      wait for delay;
      assert data_out = x"52525252525252525252525252525233" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C4";
      wait for delay;
      assert data_out = x"52525252525252525252525252525288" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C5";
      wait for delay;
      assert data_out = x"52525252525252525252525252525207" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C6";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C7" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C7";
      wait for delay;
      assert data_out = x"52525252525252525252525252525231" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C8";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B1" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000C9";
      wait for delay;
      assert data_out = x"52525252525252525252525252525212" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CA";
      wait for delay;
      assert data_out = x"52525252525252525252525252525210" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CB";
      wait for delay;
      assert data_out = x"52525252525252525252525252525259" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CC";
      wait for delay;
      assert data_out = x"52525252525252525252525252525227" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CD";
      wait for delay;
      assert data_out = x"52525252525252525252525252525280" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CE";
      wait for delay;
      assert data_out = x"525252525252525252525252525252EC" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000CF";
      wait for delay;
      assert data_out = x"5252525252525252525252525252525F" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D0";
      wait for delay;
      assert data_out = x"52525252525252525252525252525260" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D1";
      wait for delay;
      assert data_out = x"52525252525252525252525252525251" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D2";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527F" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D3";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A9" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D4";
      wait for delay;
      assert data_out = x"52525252525252525252525252525219" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D5";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B5" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D6";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D7";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520D" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D8";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522D" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000D9";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E5" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DA";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DB";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529F" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DC";
      wait for delay;
      assert data_out = x"52525252525252525252525252525293" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DD";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C9" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DE";
      wait for delay;
      assert data_out = x"5252525252525252525252525252529C" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000DF";
      wait for delay;
      assert data_out = x"525252525252525252525252525252EF" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E0";
      wait for delay;
      assert data_out = x"525252525252525252525252525252A0" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E1";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E0" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E2";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523B" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E3";
      wait for delay;
      assert data_out = x"5252525252525252525252525252524D" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E4";
      wait for delay;
      assert data_out = x"525252525252525252525252525252AE" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E5";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522A" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E6";
      wait for delay;
      assert data_out = x"525252525252525252525252525252F5" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E7";
      wait for delay;
      assert data_out = x"525252525252525252525252525252B0" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E8";
      wait for delay;
      assert data_out = x"525252525252525252525252525252C8" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000E9";
      wait for delay;
      assert data_out = x"525252525252525252525252525252EB" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000EA";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BB" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000EB";
      wait for delay;
      assert data_out = x"5252525252525252525252525252523C" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000EC";
      wait for delay;
      assert data_out = x"52525252525252525252525252525283" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000ED";
      wait for delay;
      assert data_out = x"52525252525252525252525252525253" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000EE";
      wait for delay;
      assert data_out = x"52525252525252525252525252525299" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000EF";
      wait for delay;
      assert data_out = x"52525252525252525252525252525261" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F0";
      wait for delay;
      assert data_out = x"52525252525252525252525252525217" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F1";
      wait for delay;
      assert data_out = x"5252525252525252525252525252522B" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F2";
      wait for delay;
      assert data_out = x"52525252525252525252525252525204" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F3";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527E" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F4";
      wait for delay;
      assert data_out = x"525252525252525252525252525252BA" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F5";
      wait for delay;
      assert data_out = x"52525252525252525252525252525277" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F6";
      wait for delay;
      assert data_out = x"525252525252525252525252525252D6" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F7";
      wait for delay;
      assert data_out = x"52525252525252525252525252525226" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F8";
      wait for delay;
      assert data_out = x"525252525252525252525252525252E1" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000F9";
      wait for delay;
      assert data_out = x"52525252525252525252525252525269" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FA";
      wait for delay;
      assert data_out = x"52525252525252525252525252525214" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FB";
      wait for delay;
      assert data_out = x"52525252525252525252525252525263" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FC";
      wait for delay;
      assert data_out = x"52525252525252525252525252525255" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FD";
      wait for delay;
      assert data_out = x"52525252525252525252525252525221" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FE";
      wait for delay;
      assert data_out = x"5252525252525252525252525252520C" report "Inverse SBox wrong" severity error;
      data_in <= x"000000000000000000000000000000FF";
      wait for delay;
      assert data_out = x"5252525252525252525252525252527D" report "Inverse SBox wrong" severity error;
   end process;
end ISBoxTb;